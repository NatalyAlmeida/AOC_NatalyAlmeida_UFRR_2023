library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity and1 is
    Port ( 
           entrada_a, entrada_b: in STD_LOGIC_VECTOR (15 downto 0);
           saidaComp  : out STD_LOGIC_VECTOR (15 downto 0));
end and1;

architecture andlogic of and1 is
begin
	saidaComp <= 	entrada_a AND entrada_b;
end andlogic;
